module showtime(   
    input clk,
    input reset, 
    input reg_N,
    input [6:0] wait_time,  // �ȴ�ʱ�䣨��ʱδʹ�ã�
    input [4:0] hours,      // ��ǰСʱ (Ĭ��ֵ)
    input [5:0] minutes,    // ��ǰ���� (Ĭ��ֵ)
    input [5:0] seconds,    // ��ǰ���� (Ĭ��ֵ)
    input [6:0] work_limit, // ����ʱ�����ƣ���ʱδʹ�ã�
    input power_state, 
    input [3:0] mode_state, // ģʽ״̬����ʱδʹ�ã�
    input down,             // �����¼������ڲ�ѯģʽ���л���ʾ
    output reg [3:0] an,    // Ƭѡ�ź�
    output reg [3:0] an2,   // �ڶ���Ƭѡ�ź�
    output reg [7:0] sseg,  // ��ѡ�ź�
    output reg [7:0] sseg2  // �ڶ����ѡ�ź�
);
    localparam  OFF = 1'b0,
                ON = 1'b1,
                WAITING = 1'b0,
                WORKING = 1'b1,
                MUNU = 4'b0000,
                LOW_GEAR = 4'b0001,        // һ��ģʽ
                MID_GEAR = 4'b0010,        // ����ģʽ
                HIGH_GEAR = 4'b0011,       // ����ģʽ
                AUTO_CLEAN = 4'b0100,      // �Զ����ģʽ
                MANUAL_CLEAN = 4'b0101,    // �ֶ����ģʽ
                QUERY = 4'b0110,           // ��ѯģʽ
                SET_CURRENT_TIME = 4'b0111,// ���õ�ǰʱ��ģʽ
                SET_REMINDER_TIME = 4'b1000, // ��������ʱ��ģʽ
                SET_GESTURE_TIME = 4'b1001;  // ��������ʱ��ģʽ

    // �� hex ��ֵ����Сʱ�����ӡ����Ӳ��Ϊ��λ��ʮλ����
    wire [3:0] hex0, hex1, hex2, hex3, hex4, hex5, hex6, hex7;
    
    // ��ʱ�䰴λ�ָ�Ϊʮλ�͸�λ��������ʾ���������
    assign hex0 = seconds % 10;      // ���Ӹ�λ
    assign hex1 = seconds / 10;      // ����ʮλ
    assign hex2 = minutes % 10;      // ���Ӹ�λ
    assign hex3 = minutes / 10;      // ����ʮλ
    assign hex4 = hours % 10;        // Сʱ��λ
    assign hex5 = hours / 10;        // Сʱʮλ

    localparam N = 18; // ʱ�ӷ�Ƶϵ��
    reg [3:0] hex_in, hex_in2; // ����ѡ����ʾ������
    reg [3:0] hex6_in, hex7_in; // ����ѡ����ʾhex6��hex7������
    
    // ����ģʽ״̬����hex6��hex7����ʾ
    always@* begin
        if (power_state == ON) begin // ����power_stateΪONʱ�ſ�����ʾ
            case(mode_state)
                SET_REMINDER_TIME: begin
                    hex6_in = work_limit % 10;
                    hex7_in = work_limit / 10;
                end
                SET_GESTURE_TIME: begin
                    hex6_in = wait_time % 10;
                    hex7_in = wait_time / 10;
                end
                QUERY: begin
                    if(down) begin
                        hex6_in = wait_time % 10;
                        hex7_in = wait_time / 10;
                    end else begin
                        hex6_in = work_limit % 10;
                        hex7_in = work_limit / 10;
                    end
                end
                default: begin
                    hex6_in = 4'b1111;
                    hex7_in = 4'b1111;
                end
            endcase
        end else begin
            hex6_in = 4'b1111; // power_stateΪOFFʱ����ʾ
            hex7_in = 4'b1111; // power_stateΪOFFʱ����ʾ
        end
    end
    
    // ���Ƶ�һ������ܣ���ʾ���Ӻͷ��ӣ�
    always@* begin
        if (power_state == ON) begin // ����power_stateΪONʱ�Ÿ�����ʾ
            case(regN[N-1:N-2])
                2'b00: begin
                    an = 4'b1110; // ѡ�е�1�������
                    hex_in = hex0; // ��ʾ���Ӹ�λ
                end
                2'b01: begin
                    an = 4'b1101; // ѡ�еڶ��������
                    hex_in = hex1; // ��ʾ����ʮλ
                end
                2'b10: begin
                    an = 4'b1011; // ѡ�е����������
                    hex_in = hex2; // ��ʾ���Ӹ�λ
                end
                default: begin
                    an = 4'b0111; // ѡ�е��ĸ������
                    hex_in = hex3; // ��ʾ����ʮλ
                end
            endcase
        end else begin
            an = 4'b1111; // power_stateΪOFFʱ����ʾ
            hex_in = 4'b1111; // power_stateΪOFFʱ����ʾ
        end
    end
    
    // ���Ƶڶ�������ܣ���ʾСʱ�͹���ʱ�䣩
    always@* begin
        if (power_state == ON) begin // ����power_stateΪONʱ�Ÿ�����ʾ
            case(regN[N-1:N-2])
                2'b00: begin
                    an2 = 4'b1110; // ѡ�е�1�������
                    hex_in2 = hex4; // ��ʾСʱ��λ
                end
                2'b01: begin
                    an2 = 4'b1101; // ѡ�еڶ��������
                    hex_in2 = hex5; // ��ʾСʱʮλ
                end
                2'b10: begin
                    an2 = 4'b1011; // ѡ�е����������
                    hex_in2 = hex6_in; // ��ʾ��������ʱ�������ʱ��ĸ�λ
                end
                2'b11: begin
                    an2 = 4'b0111; // ѡ�е��ĸ������
                    hex_in2 = hex7_in; // ��ʾ��������ʱ�������ʱ���ʮλ
                end
                default: begin
                    an2 = 4'b1111; // ����ʾ
                    hex_in2 = 4'b1111; // ����ʾ
                end
            endcase
        end else begin
            an2 = 4'b1111; // power_stateΪOFFʱ����ʾ
            hex_in2 = 4'b1111; // power_stateΪOFFʱ����ʾ
        end
    end
    
    // ���Ƶ�һ������������ʾ
    always@* begin
        if (power_state == ON) begin // ����power_stateΪONʱ�Ÿ�����ʾ
            case(hex_in)
                4'h0: sseg[6:0] = 7'b0000001; // ��ʾ 0
                4'h1: sseg[6:0] = 7'b1001111; // ��ʾ 1
                4'h2: sseg[6:0] = 7'b0010010; // ��ʾ 2
                4'h3: sseg[6:0] = 7'b0000110; // ��ʾ 3
                4'h4: sseg[6:0] = 7'b1001100; // ��ʾ 4
                4'h5: sseg[6:0] = 7'b0100100; // ��ʾ 5
                4'h6: sseg[6:0] = 7'b0100000; // ��ʾ 6
                4'h7: sseg[6:0] = 7'b0001111; // ��ʾ 7
                4'h8: sseg[6:0] = 7'b0000010; // ��ʾ 8
                4'h9: sseg[6:0] = 7'b0000100; // ��ʾ 9
                default: sseg[6:0] = 7'b0111000; // ��ʾĬ��ֵ
            endcase
        end else begin
            sseg[6:0] = 7'b1111111; // power_stateΪOFFʱ����ʾ
        end
    end
    
    // ���Ƶڶ�������������ʾ
    always@* begin
        if (power_state == ON) begin // ����power_stateΪONʱ�Ÿ�����ʾ
            case(hex_in2)
                4'h0: sseg2[6:0] = 7'b0000001; // ��ʾ 0
                4'h1: sseg2[6:0] = 7'b1001111; // ��ʾ 1
                4'h2: sseg2[6:0] = 7'b0010010; // ��ʾ 2
                4'h3: sseg2[6:0] = 7'b0000110; // ��ʾ 3
                4'h4: sseg2[6:0] = 7'b1001100; // ��ʾ 4
                4'h5: sseg2[6:0] = 7'b0100100; // ��ʾ 5
                4'h6: sseg2[6:0] = 7'b0100000; // ��ʾ 6
                4'h7: sseg2[6:0] = 7'b0001111; // ��ʾ 7
                4'h8: sseg2[6:0] = 7'b0000010; // ��ʾ 8
                4'h9: sseg2[6:0] = 7'b0000100; // ��ʾ 9
                default: sseg2[6:0] = 7'b0111000; // ��ʾĬ��ֵ
            endcase
        end else begin
            sseg2[6:0] = 7'b1111111; // power_stateΪOFFʱ����ʾ
        end
    end

endmodule
